/*
 * Copyright (c) 2025 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

// Change the name of this module to something that reflects its functionality and includes your name for uniqueness
// For example tqvp_yourname_spi for an SPI peripheral.
// Then edit tt_wrapper.v line 41 and change tqvp_example to your chosen module name.
module tqv_video_controller (
    input         clk,          // Clock - the TinyQV project clock is normally set to 64MHz.
    input         rst_n,        // Reset_n - low to reset.

    input  [7:0]  ui_in,        // The input PMOD, always available.  Note that ui_in[7] is normally used for UART RX.
                                // The inputs are synchronized to the clock, note this will introduce 2 cycles of delay on the inputs.

    output [7:0]  uo_out,       // The output PMOD.  Each wire is only connected if this peripheral is selected.
                                // Note that uo_out[0] is normally used for UART TX.

    input [5:0]   address,      // Address within this peripheral's address space
    input [31:0]  data_in,      // Data in to the peripheral, bottom 8, 16 or all 32 bits are valid on write.

    // Data read and write requests from the TinyQV core.
    input [1:0]   data_write_n, // 11 = no write, 00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    input [1:0]   data_read_n,  // 11 = no read,  00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    
    output [31:0] data_out,     // Data out from the peripheral, bottom 8, 16 or all 32 bits are valid on read when data_ready is high.
    output        data_ready,

    output        user_interrupt  // Dedicated interrupt request for this peripheral
);

    // Implement a 32-bit read/write register at address 0
    reg [31:0] control_data;
    always @(posedge clk) begin
        if (!rst_n) begin
            control_data <= 0;
        end else begin
            if (address == 6'h0) begin
                if (data_write_n != 2'b11)              control_data[7:0]   <= data_in[7:0];
                if (data_write_n[1] != data_write_n[0]) control_data[15:8]  <= data_in[15:8];
                if (data_write_n == 2'b10)              control_data[31:16] <= data_in[31:16];
            end
        end
    end

    // The bottom 8 bits of the stored data are added to ui_in and output to uo_out.
    //assign uo_out = example_data[7:0] + ui_in;

    wire hsync, vsync ,display_on;
    wire [9:0] hpos, ypos ;
    
    
    video_controller inst (
        .clk (clk),
        .rst (rst),
        .hsync (hsync),
        .vsync (vsync),
        .display_on(display_on),
        .hpos (hpos),
        .ypos (ypos)
    );

    reg [15:0] pix_x ;
    reg [15:0] pix_y ;

    always @ (posedge clk ) begin
        if (~rst) begin
            pix_x <= 0;
            pix_y <= 0;
        end
        else begin
            pix_x = {6'b0,hpos} ;
            pix_y = {6'b0, ypos} ;
        end
    
    end
    // Address 0 reads the example data register.  
    // Address 4 reads ui_in
    // All other addresses read 0.
    assign data_out = (address == 6'h0) ? control_data :
        (address == 6'h4) ? {16'b0, pix_x}:
        (address == 6'h6) ? {16'h0, pix_y} :
                      32'h0;

    assign uo_out[2] = hsync ;
    assign uo_out[3] = vsync ;
    assign uo_out[4] = display_on ;

    // All reads complete in 1 clock
    assign data_ready = 1;
    
    // User interrupt is generated on rising edge of ui_in[6], and cleared by writing a 1 to the low bit of address 8.
    reg example_interrupt;
    reg last_ui_in_6;

    always @(posedge clk) begin
        if (!rst_n) begin
            example_interrupt <= 0;
        end

        if (ui_in[6] && !last_ui_in_6) begin
            example_interrupt <= 1;
        end else if (address == 6'h8 && data_write_n != 2'b11 && data_in[0]) begin
            example_interrupt <= 0;
        end

        last_ui_in_6 <= ui_in[6];
    end

    assign user_interrupt = example_interrupt;

    // List all unused inputs to prevent warnings
    // data_read_n is unused as none of our behaviour depends on whether
    // registers are being read.
    wire _unused = &{data_read_n, 1'b0};

endmodule
